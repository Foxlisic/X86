module seg7
(
    input        c,
    input        e,     // =1 Активировать
    input  [3:0] d4,
    output [6:0] hex
);

reg [13:0] k; always @(posedge c) k <= k + 1;

assign hex = (e == 0) || k[13:12] ? 7'h7F : (
    //                6543210
    d4 == 4'b0000 ? 7'b1000000 : // 0
    d4 == 4'b0001 ? 7'b1111001 : // 1
    d4 == 4'b0010 ? 7'b0100100 : // 2
    d4 == 4'b0011 ? 7'b0110000 : // 3
    d4 == 4'b0100 ? 7'b0011001 : // 4
    d4 == 4'b0101 ? 7'b0010010 : // 5
    d4 == 4'b0110 ? 7'b0000010 : // 6
    d4 == 4'b0111 ? 7'b1111000 : // 7
    d4 == 4'b1000 ? 7'b0000000 : // 8
    d4 == 4'b1001 ? 7'b0010000 : // 9
    d4 == 4'b1010 ? 7'b0001000 : // A
    d4 == 4'b1011 ? 7'b0000011 : // B
    d4 == 4'b1100 ? 7'b1000110 : // C
    d4 == 4'b1101 ? 7'b0100001 : // D
    d4 == 4'b1110 ? 7'b0000110 : // E
                    7'b0001110); // F

endmodule
